magic
tech scmos
timestamp 1653039801
<< polysilicon >>
rect 12 92 15 94
rect 12 12 15 88
rect 12 5 15 8
<< ndiffusion >>
rect 8 8 12 12
rect 15 8 20 12
<< pdiffusion >>
rect 8 88 12 92
rect 15 88 20 92
<< metal1 >>
rect 4 92 8 96
rect 20 12 24 88
rect 4 4 8 8
<< metal2 >>
rect 0 96 4 100
rect 8 96 28 100
rect 0 0 4 4
rect 8 0 28 4
<< ntransistor >>
rect 12 8 15 12
<< ptransistor >>
rect 12 88 15 92
<< ndcontact >>
rect 4 8 8 12
rect 20 8 24 12
<< pdcontact >>
rect 4 88 8 92
rect 20 88 24 92
<< m2contact >>
rect 4 96 8 100
rect 4 0 8 4
<< end >>
