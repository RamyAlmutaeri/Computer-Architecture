magic
tech scmos
timestamp 1653419601
<< metal1 >>
rect 760 276 1324 280
rect 892 268 1308 272
rect 1332 200 1351 203
rect 744 188 748 199
rect 1280 188 1284 200
rect 1868 188 1872 199
rect 2404 188 2432 192
rect 264 153 268 157
rect 800 153 804 157
rect 1388 153 1392 157
rect 1924 153 1928 157
rect 204 88 220 92
rect 1328 88 1344 91
rect 180 4 184 88
rect 744 76 748 88
rect 1280 76 1284 88
rect 1868 76 1872 88
rect 2404 76 2408 80
rect 264 41 268 45
rect 800 41 804 45
rect 1388 41 1392 45
rect 1924 41 1928 45
rect 2428 4 2432 188
rect 180 0 2432 4
<< metal2 >>
rect 1312 268 1488 272
rect 888 260 1480 264
rect 880 252 1468 256
rect 1295 236 1344 240
rect 224 200 264 203
rect 224 132 228 200
rect 748 199 800 203
rect 1284 200 1328 203
rect 1355 199 1384 203
rect 1872 200 1921 203
rect 184 88 200 92
rect 224 88 264 91
rect 748 88 800 91
rect 1284 88 1324 91
rect 1348 88 1388 91
rect 1872 88 1924 91
rect 1296 20 1345 24
<< m2contact >>
rect 1308 268 1312 272
rect 884 260 888 264
rect 876 252 880 256
rect 1468 252 1472 256
rect 264 199 268 203
rect 744 199 748 203
rect 800 199 804 203
rect 1280 200 1284 204
rect 1328 200 1332 204
rect 1351 199 1355 203
rect 1384 199 1388 203
rect 1868 199 1872 203
rect 1921 200 1925 204
rect 180 88 184 92
rect 200 88 204 92
rect 220 88 224 92
rect 264 88 268 92
rect 744 88 748 92
rect 800 88 804 92
rect 1280 88 1284 92
rect 1324 88 1328 92
rect 1344 88 1348 92
rect 1388 88 1392 92
rect 1868 88 1872 92
rect 1924 88 1928 92
use 4in-multiplier  4in-multiplier_0
timestamp 1653191793
transform 1 0 900 0 1 132
box -708 -120 400 148
use 4in-multiplier  4in-multiplier_1
timestamp 1653191793
transform 1 0 2024 0 1 132
box -708 -120 400 148
<< end >>
