magic
tech scmos
timestamp 1653420455
<< error_s >>
rect 1747 2372 1751 2374
rect 2875 2372 2879 2374
rect 4003 2372 4007 2374
rect 10208 1443 10214 1446
<< metal1 >>
rect -92 2764 4483 2768
rect -92 2188 -88 2764
rect -3568 2184 -88 2188
rect -80 2752 3947 2756
rect -80 2176 -76 2752
rect -2476 2172 -76 2176
rect -68 2740 3355 2744
rect -68 2164 -64 2740
rect -1360 2160 -64 2164
rect -56 2728 2819 2732
rect -56 2152 -52 2728
rect -44 2716 2227 2720
rect -44 2168 -40 2716
rect -32 2704 1690 2708
rect -32 2180 -28 2704
rect -20 2692 1098 2696
rect -20 2192 -16 2692
rect -8 2680 563 2684
rect -8 2204 -4 2680
rect 2312 2667 2316 2671
rect 2312 2655 2316 2659
rect 2312 2639 2316 2643
rect 2312 2619 2316 2623
rect 563 2567 567 2611
rect 571 2524 575 2611
rect 1099 2567 1103 2611
rect 1108 2524 1111 2611
rect 1691 2567 1694 2612
rect 1699 2524 1702 2611
rect 2227 2567 2231 2611
rect 2239 2524 2243 2611
rect 2819 2567 2823 2611
rect 2827 2524 2830 2612
rect 3355 2569 3359 2612
rect 3368 2612 3369 2613
rect 3364 2524 3369 2612
rect 3947 2567 3951 2611
rect 3956 2524 3959 2611
rect 4483 2555 4487 2611
rect 24 2520 45 2523
rect 1153 2520 1174 2524
rect 2280 2520 2300 2524
rect 3364 2520 3365 2524
rect 3412 2520 3428 2524
rect 23 2408 48 2411
rect 563 2383 566 2448
rect 619 2373 623 2412
rect 1099 2380 1103 2447
rect 1211 2380 1215 2412
rect 1691 2380 1695 2447
rect 1747 2376 1751 2412
rect 2227 2380 2231 2446
rect 2339 2380 2343 2412
rect 2818 2383 2823 2446
rect 2818 2380 2819 2383
rect 2875 2376 2879 2408
rect 3354 2383 3359 2445
rect 3467 2381 3470 2409
rect 3947 2383 3952 2446
rect 3947 2380 3948 2383
rect 4003 2377 4007 2408
rect 4003 2372 4007 2373
rect 1060 2216 1064 2363
rect 1099 2292 1103 2328
rect 1691 2297 1695 2323
rect 2227 2296 2231 2324
rect 2819 2316 2824 2317
rect 2819 2296 2824 2312
rect 3354 2292 3358 2322
rect 3947 2317 3948 2320
rect 3947 2295 3952 2317
rect 1099 2284 1104 2292
rect 3947 2291 3948 2295
rect 1099 2280 11796 2284
rect 1695 2268 10704 2272
rect 2231 2256 9620 2260
rect 2824 2245 8524 2249
rect 3359 2236 7412 2240
rect 3951 2224 6292 2227
rect 3947 2223 6292 2224
rect 1060 2212 5223 2216
rect -8 2200 4108 2204
rect -20 2188 3024 2192
rect -32 2176 1896 2180
rect -44 2164 812 2168
rect -292 2148 -52 2152
rect 13395 1551 17844 1556
rect -753 1443 -748 1447
rect 331 1443 336 1447
rect 1431 1443 1436 1447
rect 2515 1443 2520 1447
rect 3631 1443 3636 1447
rect 4715 1443 4720 1447
rect 5831 1443 5836 1447
rect 6915 1443 6920 1447
rect -3488 1383 -3484 1431
rect -3488 908 -3484 1332
rect -2957 924 -2953 1443
rect -2404 1383 -2400 1431
rect -2404 1336 -2400 1340
rect -2404 920 -2400 1332
rect -1873 932 -1869 1443
rect -1292 1383 -1287 1431
rect -1288 1381 -1287 1383
rect -1292 932 -1288 1340
rect -752 940 -748 1443
rect -207 1383 -203 1431
rect -207 1336 -203 1352
rect -207 944 -203 1332
rect 332 952 336 1443
rect 897 1383 900 1432
rect 896 1335 900 1345
rect 896 956 900 1331
rect 1432 964 1436 1443
rect 1984 1383 1987 1431
rect 1984 1336 1988 1343
rect 1984 968 1988 1332
rect 2516 976 2520 1443
rect 3092 1383 3097 1430
rect 3096 1380 3097 1383
rect 3092 1336 3096 1344
rect 3092 980 3096 1332
rect 3092 976 3484 980
rect 1984 964 2872 968
rect 896 952 2344 956
rect -207 940 1752 944
rect -1292 928 1268 932
rect -2404 916 616 920
rect -3488 904 216 908
rect -2957 153 -2953 896
rect -1873 320 -1869 896
rect -752 392 -748 896
rect -752 388 -116 392
rect -1873 316 -112 320
rect -2957 149 -108 153
rect -100 -79 -96 708
rect -88 -68 -84 692
rect -76 -56 -72 680
rect -64 -44 -60 668
rect -52 -32 -48 652
rect -40 -20 -36 640
rect -28 -8 -24 628
rect -12 12 -8 616
rect 4 388 200 392
rect 124 368 204 372
rect 124 288 128 368
rect 212 296 216 904
rect 228 388 320 392
rect 332 380 336 908
rect 563 708 564 712
rect 568 708 628 712
rect 580 692 642 696
rect 600 680 628 684
rect 588 668 632 672
rect 608 652 632 656
rect 608 640 632 644
rect 608 628 632 632
rect 608 616 632 620
rect 348 388 1156 392
rect 224 368 1248 372
rect 332 308 336 360
rect 540 356 1248 360
rect 332 304 532 308
rect 540 288 544 356
rect 552 304 1240 308
rect 1248 288 1252 344
rect 1264 296 1268 928
rect 1432 384 1436 932
rect 1728 708 1729 712
rect 1733 708 1765 712
rect 1741 692 1742 696
rect 1746 692 1765 696
rect 1740 680 1761 684
rect 1728 668 1764 672
rect 1736 652 1764 656
rect 1744 640 1764 644
rect 1744 628 1764 632
rect 1744 616 1764 620
rect 1432 380 2288 384
rect 1280 368 2328 372
rect 1280 356 2328 360
rect 1280 344 2328 348
rect 1664 332 2328 336
rect 1276 304 1652 308
rect 1664 288 1668 332
rect 1684 284 1688 304
rect 2340 296 2344 952
rect 2516 384 2520 956
rect 2844 708 2884 712
rect 2844 692 2884 696
rect 2848 680 2884 684
rect 2860 668 2884 672
rect 2868 652 2884 656
rect 2860 640 2884 644
rect 2860 628 2884 632
rect 2860 616 2884 620
rect 2516 380 2808 384
rect 3408 376 3468 380
rect 2356 368 3468 372
rect 2356 356 3468 360
rect 2356 344 3468 348
rect 2356 332 3468 336
rect 2372 320 3468 324
rect 2372 288 2376 320
rect 2788 304 3468 308
rect 2788 284 2792 304
rect 3480 296 3484 976
rect 3632 380 3636 1443
rect 4183 1383 4186 1431
rect 4183 996 4187 1342
rect 3988 992 4187 996
rect 4716 720 4720 1443
rect 5301 1383 5304 1430
rect 3952 708 5284 712
rect 3952 692 5284 696
rect 3960 680 5288 684
rect 3968 668 5288 672
rect 3976 652 5272 656
rect 3980 640 5284 644
rect 3980 628 5284 632
rect 5301 620 5305 1363
rect 5832 720 5836 1443
rect 6384 1383 6387 1431
rect 5316 708 6348 712
rect 5316 692 6348 696
rect 5320 680 6360 684
rect 5320 668 6368 672
rect 5316 652 6368 656
rect 5316 640 6376 644
rect 6384 632 6388 1358
rect 6916 728 6920 1443
rect 7500 1383 7504 1431
rect 6396 708 7456 712
rect 6396 692 7456 696
rect 6396 680 7464 684
rect 6396 668 7472 672
rect 6396 652 7448 656
rect 7500 644 7504 1361
rect 8027 724 8031 1443
rect 8583 1383 8588 1430
rect 8587 1380 8588 1383
rect 7512 708 8557 712
rect 7512 692 8556 696
rect 7516 680 8568 684
rect 7516 668 8575 672
rect 8584 656 8588 1357
rect 9111 728 9115 1443
rect 9681 1383 9685 1431
rect 8598 708 9657 712
rect 8596 692 9655 696
rect 8601 680 9668 684
rect 9681 672 9685 1358
rect 10207 728 10211 1443
rect 10764 1383 10767 1431
rect 9696 708 10752 712
rect 9696 692 10752 696
rect 10764 684 10768 1360
rect 11295 728 11299 1447
rect 11876 1383 11880 1431
rect 10795 708 10796 712
rect 10800 708 11864 712
rect 11876 696 11880 1352
rect 12411 728 12415 1447
rect 13499 1443 13521 1447
rect 12964 1383 12968 1431
rect 12964 712 12968 1352
rect 11888 708 12968 712
rect 10800 692 11880 696
rect 9696 680 10768 684
rect 8600 668 9685 672
rect 7516 652 8588 656
rect 6392 640 6393 644
rect 6397 640 7504 644
rect 5316 628 6388 632
rect 3980 616 5305 620
rect 3496 376 3636 380
rect 4712 380 4716 608
rect 5832 372 5836 620
rect 3496 368 5836 372
rect 6916 360 6920 632
rect 3496 356 6920 360
rect 8027 348 8031 640
rect 3496 344 8031 348
rect 9111 336 9116 652
rect 3496 332 9116 336
rect 10207 324 10211 668
rect 3496 320 10211 324
rect 3496 304 11295 308
rect 12411 300 12415 684
rect 3516 296 12415 300
rect 3516 288 3520 296
rect 4712 284 4716 288
rect 3936 280 4716 284
rect 3912 272 3916 276
rect 13518 268 13521 1443
rect 17244 993 17248 997
rect 17244 985 17248 989
rect 17244 977 17248 981
rect 17244 969 17248 973
rect 16153 874 16156 961
rect 17278 874 17281 961
rect 17892 956 17896 2604
rect 17828 952 17896 956
rect 15610 870 15636 874
rect 15640 870 15641 874
rect 16737 870 16752 874
rect 15606 757 15620 761
rect 15624 757 15625 761
rect 16202 731 16206 761
rect 16699 732 16702 870
rect 16730 758 16745 762
rect 16707 732 16710 758
rect 17326 731 17329 762
rect 3912 264 3916 268
rect 4080 264 13521 268
rect 124 228 128 264
rect 3912 256 3916 260
rect 3912 248 3916 252
rect 16 149 72 153
rect 124 116 128 140
rect 540 41 544 240
rect 560 228 564 240
rect 1156 228 1160 240
rect 1248 228 1252 240
rect 552 186 556 189
rect 1088 186 1092 189
rect 1248 112 1252 140
rect 1088 61 1092 64
rect 552 57 556 60
rect 1664 41 1668 240
rect 1684 228 1688 240
rect 1676 186 1680 189
rect 2212 186 2216 189
rect 2236 153 2240 240
rect 2372 228 2376 240
rect 2372 116 2376 140
rect 1676 66 1680 69
rect 2212 68 2216 71
rect 2788 41 2792 240
rect 2808 228 2812 240
rect 3404 224 3408 240
rect 2800 188 2804 191
rect 3336 188 3340 191
rect 2800 61 2804 64
rect 3336 52 3340 55
rect 72 24 76 37
rect 124 24 128 28
rect 72 20 128 24
rect 1196 24 1200 37
rect 1196 20 1252 24
rect 2320 24 2324 41
rect 2372 24 2376 28
rect 3444 28 3448 37
rect 3516 28 3520 240
rect 3932 228 3936 240
rect 4080 228 4084 264
rect 17892 237 17896 952
rect 17908 740 17912 2388
rect 3924 192 3928 195
rect 4460 193 4464 196
rect 4032 112 4036 136
rect 4460 55 4464 58
rect 3924 51 3928 54
rect 3980 24 3984 37
rect 2320 20 2376 24
rect 3980 20 4036 24
rect 17908 20 17912 736
rect 588 -8 592 8
rect -28 -12 592 -8
rect -40 -24 1152 -20
rect 1720 -32 1724 12
rect -52 -36 1724 -32
rect -64 -48 2276 -44
rect -64 -49 -60 -48
rect 2836 -56 2840 12
rect -76 -60 2840 -56
rect -88 -72 3400 -68
rect 3960 -79 3964 12
rect -100 -83 3964 -79
<< metal2 >>
rect 4482 2764 4483 2768
rect 4487 2764 4488 2768
rect 3951 2752 3952 2756
rect 563 2615 567 2680
rect 571 2615 575 2684
rect 1099 2615 1103 2692
rect 1108 2615 1111 2696
rect 1690 2616 1694 2704
rect 1690 2612 1691 2616
rect 1699 2615 1702 2702
rect 2227 2615 2231 2716
rect 2239 2704 2243 2705
rect 2239 2615 2243 2700
rect 2819 2615 2823 2728
rect 2827 2616 2830 2704
rect 3355 2616 3359 2740
rect 3364 2701 3365 2705
rect 3364 2616 3369 2701
rect 3368 2612 3369 2616
rect 3947 2689 3952 2752
rect 3947 2615 3951 2689
rect 3956 2615 3959 2700
rect 4482 2667 4488 2764
rect 4483 2615 4487 2667
rect 4500 2604 17892 2607
rect 4500 2603 17896 2604
rect -98 2520 20 2523
rect 49 2520 83 2523
rect 575 2520 619 2523
rect 1112 2520 1149 2524
rect 1178 2520 1211 2524
rect 1703 2520 1747 2523
rect 2243 2520 2276 2524
rect 2280 2520 2281 2524
rect 2304 2520 2339 2524
rect 2831 2520 2875 2523
rect 3369 2520 3408 2524
rect 3432 2520 3467 2524
rect 3960 2520 4003 2523
rect -96 2408 19 2411
rect 52 2408 83 2411
rect 4499 2388 17908 2391
rect 4499 2387 17912 2388
rect 563 2308 566 2379
rect 619 2334 623 2369
rect 1099 2332 1103 2376
rect 1211 2348 1215 2376
rect 1691 2328 1695 2376
rect 1747 2340 1751 2372
rect 2227 2320 2231 2376
rect 2339 2346 2343 2376
rect 2823 2379 2824 2382
rect 2819 2316 2824 2379
rect 2875 2343 2879 2372
rect 3354 2326 3357 2379
rect 3947 2379 3948 2382
rect 3467 2351 3470 2377
rect 3947 2321 3952 2379
rect 4003 2344 4007 2373
rect 3947 2317 3948 2321
rect 3947 2316 3952 2317
rect 12912 2309 12916 2310
rect 4649 2308 12916 2309
rect 563 2304 12916 2308
rect 563 2303 4652 2304
rect 1691 2273 1695 2292
rect 2227 2260 2231 2292
rect 2819 2249 2824 2292
rect 2819 2244 2824 2245
rect 3947 2291 3948 2293
rect 3354 2240 3357 2288
rect 3947 2228 3952 2291
rect 3951 2227 3952 2228
rect -3572 1503 -3568 2184
rect -2480 1503 -2476 2172
rect -1364 1503 -1360 2160
rect -292 1504 -288 2152
rect -292 1499 -288 1500
rect 812 1503 816 2164
rect 1896 1503 1900 2176
rect 3024 1503 3028 2188
rect 4108 1503 4112 2200
rect 5223 1503 5227 2212
rect 6292 1503 6296 2222
rect 7412 1503 7416 2236
rect 8524 1503 8528 2245
rect 9620 1503 9624 2256
rect 10704 1503 10708 2268
rect 11796 1503 11800 2280
rect 12912 1503 12916 2304
rect -3488 1336 -3484 1379
rect -2404 1336 -2400 1379
rect -1292 1344 -1288 1379
rect -207 1336 -203 1379
rect 897 1335 900 1379
rect 3096 1379 3097 1383
rect 1984 1336 1987 1379
rect 3092 1336 3097 1379
rect 4183 1346 4186 1379
rect 5301 1367 5304 1379
rect 6384 1362 6387 1379
rect 8587 1379 8588 1382
rect 7500 1365 7503 1379
rect 8583 1361 8588 1379
rect 8583 1357 8584 1361
rect 9681 1362 9685 1379
rect 10764 1364 10767 1379
rect 11876 1356 11880 1379
rect 12964 1356 12968 1379
rect 3096 1333 3097 1336
rect -2957 900 -2953 920
rect -1873 900 -1869 928
rect -752 900 -748 936
rect 332 912 336 948
rect 1432 936 1436 960
rect 2516 960 2520 972
rect -96 708 564 712
rect -84 692 576 696
rect -72 680 596 684
rect -60 668 584 672
rect -48 652 604 656
rect -36 640 604 644
rect -24 628 604 632
rect -8 616 604 620
rect -112 388 0 392
rect 204 388 224 392
rect 324 388 344 392
rect 208 368 220 372
rect 332 364 336 376
rect -108 316 564 320
rect 536 304 548 308
rect 124 268 128 284
rect 540 244 544 284
rect 560 244 564 316
rect 616 244 620 916
rect 632 708 1729 712
rect 646 692 1742 696
rect 632 680 1736 684
rect 636 668 1724 672
rect 636 652 1732 656
rect 636 640 1740 644
rect 636 628 1740 632
rect 636 616 1740 620
rect 1156 244 1160 388
rect 1252 368 1276 372
rect 1252 356 1276 360
rect 1252 344 1276 348
rect 1244 304 1272 308
rect 1656 304 1684 308
rect 1248 244 1252 284
rect 1664 244 1668 284
rect 1684 244 1688 280
rect 1752 244 1756 940
rect 1769 708 2840 712
rect 1769 692 2840 696
rect 1765 680 2844 684
rect 2848 680 2849 684
rect 1768 668 2856 672
rect 1768 652 2864 656
rect 1768 640 2856 644
rect 1768 628 2856 632
rect 1768 616 2856 620
rect 2288 244 2292 380
rect 2332 368 2352 372
rect 2332 356 2352 360
rect 2332 344 2352 348
rect 2332 332 2352 336
rect 2240 240 2292 244
rect 2372 244 2376 284
rect 2788 244 2792 280
rect 2808 244 2812 380
rect 2872 244 2876 964
rect 2888 708 3948 712
rect 2888 692 3948 696
rect 2888 680 3956 684
rect 2888 668 3964 672
rect 2888 652 3972 656
rect 2888 640 3976 644
rect 2888 628 3976 632
rect 2888 616 3976 620
rect 3472 376 3492 380
rect 3404 244 3408 376
rect 3472 368 3492 372
rect 3472 356 3492 360
rect 3472 344 3492 348
rect 3472 332 3492 336
rect 3472 320 3492 324
rect 3472 304 3492 308
rect 3516 244 3520 284
rect 3932 244 3936 280
rect 3988 244 3992 995
rect 16153 965 16156 1009
rect 17278 965 17281 1036
rect 15577 870 15606 874
rect 15635 870 15636 874
rect 15640 870 15666 874
rect 16157 870 16202 874
rect 16206 870 16207 874
rect 16703 870 16733 873
rect 16756 870 16790 874
rect 17282 870 17326 873
rect 17844 796 17848 1551
rect 17810 793 17848 796
rect 15636 761 15666 762
rect 15569 757 15602 761
rect 15624 758 15666 761
rect 15670 758 15671 762
rect 16711 758 16726 762
rect 16749 758 16790 762
rect 15624 757 15655 758
rect 17823 740 17912 741
rect 17823 737 17908 740
rect 4712 612 4716 720
rect 5288 708 5312 712
rect 5288 692 5312 696
rect 5292 680 5316 684
rect 5292 668 5316 672
rect 5276 652 5312 656
rect 5288 640 5312 644
rect 5288 628 5312 632
rect 5316 628 5317 632
rect 5832 624 5836 716
rect 6352 708 6392 712
rect 6352 692 6392 696
rect 6364 680 6392 684
rect 6372 668 6392 672
rect 6372 652 6392 656
rect 6380 640 6393 644
rect 6916 636 6920 724
rect 7460 708 7508 712
rect 7460 692 7508 696
rect 7468 680 7512 684
rect 7476 668 7512 672
rect 7452 652 7512 656
rect 8027 644 8031 720
rect 8561 708 8594 712
rect 8560 692 8592 696
rect 8572 680 8597 684
rect 8579 668 8596 672
rect 9111 656 9115 724
rect 9661 708 9692 712
rect 9696 708 9698 712
rect 9659 692 9692 696
rect 9672 680 9692 684
rect 10207 672 10211 724
rect 10756 708 10796 712
rect 10756 692 10796 696
rect 4712 292 4716 376
rect 11295 308 11299 724
rect 11868 708 11884 712
rect 12411 688 12415 724
rect 16202 699 16206 727
rect 16699 704 16702 728
rect 16707 700 16710 728
rect 17326 698 17329 727
rect 4477 232 17892 236
rect -104 149 12 153
rect 124 144 128 224
rect 560 153 564 224
rect 1156 153 1160 224
rect 560 149 608 153
rect 1156 149 1196 153
rect 1248 144 1252 224
rect 1684 153 1688 224
rect 1684 149 1732 153
rect 2240 149 2320 153
rect 2372 144 2376 224
rect 2808 153 2812 224
rect 3404 153 3408 220
rect 3932 153 3936 224
rect 4032 224 4080 228
rect 2808 149 2856 153
rect 3404 149 3444 153
rect 3932 149 3976 153
rect 4032 140 4036 224
rect 124 32 128 112
rect 544 37 604 41
rect 1248 28 1252 108
rect 1668 37 1732 41
rect 2372 32 2376 112
rect 2792 37 2852 41
rect 4032 28 4036 108
rect 3448 24 3516 28
rect 4476 16 17908 20
rect -8 8 28 12
rect 1152 -20 1156 8
rect 2276 -44 2280 8
rect 3400 -68 3404 8
<< m2contact >>
rect 4483 2764 4487 2768
rect -102 2520 -98 2524
rect -100 2408 -96 2412
rect -3572 2184 -3568 2188
rect 3947 2752 3951 2756
rect -2480 2172 -2476 2176
rect 3355 2740 3359 2744
rect -1364 2160 -1360 2164
rect 2819 2728 2823 2732
rect 2227 2716 2231 2720
rect 1690 2704 1694 2708
rect 1699 2702 1703 2706
rect 2827 2704 2831 2708
rect 2239 2700 2243 2704
rect 3365 2701 3369 2705
rect 3956 2700 3960 2704
rect 1108 2696 1112 2700
rect 1098 2692 1103 2696
rect 571 2684 575 2688
rect 563 2680 567 2684
rect 563 2611 567 2615
rect 571 2611 575 2615
rect 1099 2611 1103 2615
rect 1108 2611 1112 2615
rect 1691 2612 1695 2616
rect 1699 2611 1703 2615
rect 2227 2611 2231 2615
rect 2239 2611 2243 2615
rect 2819 2611 2823 2615
rect 2827 2612 2831 2616
rect 3355 2612 3359 2616
rect 3364 2612 3368 2616
rect 3947 2611 3951 2615
rect 3955 2611 3959 2615
rect 4483 2611 4487 2615
rect 17892 2604 17896 2608
rect 20 2520 24 2524
rect 45 2520 49 2524
rect 83 2520 87 2524
rect 571 2520 575 2524
rect 619 2520 623 2524
rect 1108 2520 1112 2524
rect 1149 2520 1153 2524
rect 1174 2520 1178 2524
rect 1211 2520 1215 2524
rect 1699 2520 1703 2524
rect 1747 2520 1751 2524
rect 2239 2520 2243 2524
rect 2276 2520 2280 2524
rect 2300 2520 2304 2524
rect 2339 2520 2343 2524
rect 2827 2520 2831 2524
rect 2875 2520 2879 2524
rect 3365 2520 3369 2524
rect 3408 2520 3412 2524
rect 3428 2520 3432 2524
rect 3467 2520 3471 2524
rect 3956 2520 3960 2524
rect 4003 2520 4007 2524
rect 19 2408 23 2412
rect 48 2408 52 2412
rect 83 2408 87 2412
rect 563 2379 567 2383
rect 1099 2376 1103 2380
rect 1211 2376 1215 2380
rect 1691 2376 1695 2380
rect 2227 2376 2231 2380
rect 2339 2376 2343 2380
rect 2819 2379 2823 2383
rect 3354 2379 3359 2383
rect 3467 2377 3471 2381
rect 3948 2379 3952 2383
rect 619 2369 623 2373
rect 1747 2372 1751 2376
rect 2875 2372 2879 2376
rect 4003 2373 4007 2377
rect 619 2330 623 2334
rect 1211 2344 1215 2348
rect 3467 2347 3471 2351
rect 2339 2342 2343 2346
rect 1747 2336 1751 2340
rect 2875 2339 2879 2343
rect 4003 2340 4007 2344
rect 1099 2328 1103 2332
rect 1691 2323 1695 2328
rect 1691 2292 1695 2297
rect 3354 2322 3359 2326
rect 2227 2292 2231 2296
rect 2819 2312 2824 2316
rect 2819 2292 2824 2296
rect 3948 2317 3952 2321
rect 3354 2288 3359 2292
rect 3948 2291 3952 2295
rect 11796 2280 11800 2284
rect 1691 2268 1695 2273
rect 10704 2268 10708 2272
rect 2227 2256 2231 2260
rect 9620 2256 9624 2260
rect 2819 2245 2824 2249
rect 8524 2245 8528 2249
rect 3354 2236 3359 2240
rect 7412 2236 7416 2240
rect 3947 2224 3951 2228
rect 6292 2222 6296 2228
rect 5223 2212 5227 2216
rect 4108 2200 4112 2204
rect 3024 2188 3028 2192
rect 1896 2176 1900 2180
rect 812 2164 816 2168
rect 17844 1551 17848 1556
rect -3572 1499 -3568 1503
rect -2480 1499 -2476 1503
rect -1364 1499 -1360 1503
rect -292 1500 -288 1504
rect 812 1499 816 1503
rect 1896 1499 1900 1503
rect 3024 1499 3028 1503
rect 4108 1499 4112 1503
rect 5223 1499 5227 1503
rect 6292 1499 6296 1503
rect 7412 1499 7416 1503
rect 8524 1499 8528 1503
rect 9620 1499 9624 1503
rect 10704 1499 10708 1503
rect 11796 1499 11800 1503
rect 12912 1499 12916 1503
rect -3488 1379 -3484 1383
rect -3488 1332 -3484 1336
rect -2404 1379 -2400 1383
rect -2957 920 -2953 924
rect -2404 1332 -2400 1336
rect -1292 1379 -1288 1383
rect -1873 928 -1869 932
rect -1292 1340 -1288 1344
rect -207 1379 -203 1383
rect -207 1332 -203 1336
rect 896 1379 900 1383
rect 896 1331 900 1335
rect 1984 1379 1988 1383
rect 1984 1332 1988 1336
rect 3092 1379 3096 1383
rect 3092 1332 3096 1336
rect 2516 972 2520 976
rect 2872 964 2876 968
rect 1432 960 1436 964
rect 2516 956 2520 960
rect 332 948 336 952
rect 1752 940 1756 944
rect -752 936 -748 940
rect 1432 932 1436 936
rect 616 916 620 920
rect 332 908 336 912
rect -2957 896 -2953 900
rect -1873 896 -1869 900
rect -752 896 -748 900
rect -100 708 -96 712
rect -116 388 -112 392
rect -112 316 -108 320
rect -108 149 -104 153
rect -88 692 -84 696
rect -76 680 -72 684
rect -64 668 -60 672
rect -52 652 -48 656
rect -40 640 -36 644
rect -28 628 -24 632
rect -12 616 -8 620
rect 0 388 4 392
rect 200 388 204 392
rect 204 368 208 372
rect 224 388 228 392
rect 320 388 324 392
rect 564 708 568 712
rect 628 708 632 712
rect 576 692 580 696
rect 642 692 646 696
rect 596 680 600 684
rect 628 680 632 684
rect 584 668 588 672
rect 632 668 636 672
rect 604 652 608 656
rect 632 652 636 656
rect 604 640 608 644
rect 632 640 636 644
rect 604 628 608 632
rect 632 628 636 632
rect 604 616 608 620
rect 632 616 636 620
rect 344 388 348 392
rect 1156 388 1160 392
rect 332 376 336 380
rect 220 368 224 372
rect 1248 368 1252 372
rect 332 360 336 364
rect 1248 356 1252 360
rect 532 304 536 308
rect 212 292 216 296
rect 124 284 128 288
rect 1248 344 1252 348
rect 548 304 552 308
rect 1240 304 1244 308
rect 540 284 544 288
rect 1729 708 1733 712
rect 1765 708 1769 712
rect 1742 692 1746 696
rect 1765 692 1769 696
rect 1736 680 1740 684
rect 1761 680 1765 684
rect 1724 668 1728 672
rect 1764 668 1768 672
rect 1732 652 1736 656
rect 1764 652 1768 656
rect 1740 640 1744 644
rect 1764 640 1768 644
rect 1740 628 1744 632
rect 1764 628 1768 632
rect 1740 616 1744 620
rect 1764 616 1768 620
rect 2288 380 2292 384
rect 1276 368 1280 372
rect 2328 368 2332 372
rect 1276 356 1280 360
rect 2328 356 2332 360
rect 1276 344 1280 348
rect 2328 344 2332 348
rect 2328 332 2332 336
rect 1272 304 1276 308
rect 1652 304 1656 308
rect 1264 292 1268 296
rect 1248 284 1252 288
rect 1664 284 1668 288
rect 1684 304 1688 308
rect 2840 708 2844 712
rect 2884 708 2888 712
rect 2840 692 2844 696
rect 2884 692 2888 696
rect 2844 680 2848 684
rect 2884 680 2888 684
rect 2856 668 2860 672
rect 2884 668 2888 672
rect 2864 652 2868 656
rect 2884 652 2888 656
rect 2856 640 2860 644
rect 2884 640 2888 644
rect 2856 628 2860 632
rect 2884 628 2888 632
rect 2856 616 2860 620
rect 2884 616 2888 620
rect 2808 380 2812 384
rect 3404 376 3408 380
rect 3468 376 3472 380
rect 2352 368 2356 372
rect 3468 368 3472 372
rect 2352 356 2356 360
rect 3468 356 3472 360
rect 2352 344 2356 348
rect 3468 344 3472 348
rect 2352 332 2356 336
rect 3468 332 3472 336
rect 2340 292 2344 296
rect 3468 320 3472 324
rect 2372 284 2376 288
rect 3468 304 3472 308
rect 4182 1379 4187 1383
rect 4183 1342 4188 1346
rect 5301 1379 5305 1383
rect 4716 716 4720 720
rect 5301 1363 5305 1367
rect 3948 708 3952 712
rect 5284 708 5288 712
rect 3948 692 3952 696
rect 5284 692 5288 696
rect 3956 680 3960 684
rect 5288 680 5292 684
rect 3964 668 3968 672
rect 5288 668 5292 672
rect 3972 652 3976 656
rect 5272 652 5276 656
rect 3976 640 3980 644
rect 5284 640 5288 644
rect 3976 628 3980 632
rect 5284 628 5288 632
rect 6383 1379 6387 1383
rect 5832 716 5836 720
rect 6384 1358 6388 1362
rect 5312 708 5316 712
rect 6348 708 6352 712
rect 5312 692 5316 696
rect 6348 692 6352 696
rect 5316 680 5320 684
rect 6360 680 6364 684
rect 5316 668 5320 672
rect 6368 668 6372 672
rect 5312 652 5316 656
rect 6368 652 6372 656
rect 5312 640 5316 644
rect 6376 640 6380 644
rect 7500 1379 7504 1383
rect 6916 724 6920 728
rect 7500 1361 7504 1365
rect 6392 708 6396 712
rect 7456 708 7460 712
rect 6392 692 6396 696
rect 7456 692 7460 696
rect 6392 680 6396 684
rect 7464 680 7468 684
rect 6392 668 6396 672
rect 7472 668 7476 672
rect 6392 652 6396 656
rect 7448 652 7452 656
rect 8583 1379 8587 1383
rect 8027 720 8031 724
rect 8584 1357 8588 1361
rect 7508 708 7512 712
rect 8557 708 8561 712
rect 7508 692 7512 696
rect 8556 692 8560 696
rect 7512 680 7516 684
rect 8568 680 8572 684
rect 7512 668 7516 672
rect 8575 668 8579 672
rect 9681 1379 9685 1383
rect 9681 1358 9685 1362
rect 9111 724 9116 728
rect 8594 708 8598 712
rect 9657 708 9661 712
rect 8592 692 8596 696
rect 9655 692 9659 696
rect 8597 680 8601 684
rect 9668 680 9672 684
rect 10764 1379 10768 1383
rect 10207 724 10211 728
rect 10764 1360 10768 1364
rect 9692 708 9696 712
rect 10752 708 10756 712
rect 9692 692 9696 696
rect 10752 692 10756 696
rect 11876 1379 11880 1383
rect 11295 724 11299 728
rect 11876 1352 11880 1356
rect 10796 708 10800 712
rect 11864 708 11868 712
rect 12964 1379 12968 1383
rect 12411 724 12415 728
rect 12964 1352 12968 1356
rect 11884 708 11888 712
rect 10796 692 10800 696
rect 9692 680 9696 684
rect 12411 684 12415 688
rect 8596 668 8600 672
rect 10207 668 10211 672
rect 7512 652 7516 656
rect 9111 652 9116 656
rect 6393 640 6397 644
rect 8027 640 8031 644
rect 5312 628 5316 632
rect 6916 632 6920 636
rect 3976 616 3980 620
rect 5832 620 5836 624
rect 3492 376 3496 380
rect 4712 608 4716 612
rect 4712 376 4716 380
rect 3492 368 3496 372
rect 3492 356 3496 360
rect 3492 344 3496 348
rect 3492 332 3496 336
rect 3492 320 3496 324
rect 3492 304 3496 308
rect 11295 304 11299 308
rect 3480 292 3484 296
rect 3516 284 3520 288
rect 4712 288 4716 292
rect 1684 280 1688 284
rect 2788 280 2792 284
rect 3932 280 3936 284
rect 17278 1036 17282 1040
rect 16152 1009 16156 1013
rect 16153 961 16157 965
rect 17278 961 17282 965
rect 17824 952 17828 956
rect 15573 870 15577 874
rect 15606 870 15610 874
rect 15636 870 15640 874
rect 15666 870 15670 874
rect 16153 870 16157 874
rect 16202 870 16206 874
rect 16699 870 16703 874
rect 16733 870 16737 874
rect 16752 870 16756 874
rect 16790 870 16794 874
rect 17278 870 17282 874
rect 17326 870 17330 874
rect 15565 757 15569 761
rect 15602 757 15606 761
rect 15620 757 15624 761
rect 15666 758 15670 762
rect 16202 727 16206 731
rect 17806 793 17810 798
rect 16707 758 16711 762
rect 16726 758 16730 762
rect 16745 758 16749 762
rect 16790 758 16794 762
rect 16699 728 16703 732
rect 16707 728 16711 732
rect 17326 727 17330 731
rect 16699 700 16703 704
rect 16202 695 16206 699
rect 16707 696 16711 700
rect 17326 694 17330 698
rect 124 264 128 268
rect 124 224 128 228
rect 540 240 544 244
rect 12 149 16 153
rect 124 140 128 144
rect 124 112 128 116
rect 560 240 564 244
rect 616 240 620 244
rect 1156 240 1160 244
rect 560 224 564 228
rect 1156 224 1160 228
rect 1248 240 1252 244
rect 1248 224 1252 228
rect 1664 240 1668 244
rect 1196 149 1200 153
rect 1248 140 1252 144
rect 1248 108 1252 112
rect 1684 240 1688 244
rect 1752 240 1756 244
rect 2236 240 2240 244
rect 1684 224 1688 228
rect 2372 240 2376 244
rect 2372 224 2376 228
rect 2788 240 2792 244
rect 1732 149 1736 153
rect 2236 149 2240 153
rect 2372 140 2376 144
rect 2372 112 2376 116
rect 2808 240 2812 244
rect 2872 240 2876 244
rect 3404 240 3408 244
rect 2808 224 2812 228
rect 3404 220 3408 224
rect 3516 240 3520 244
rect 2856 149 2860 153
rect 3444 149 3448 153
rect 540 37 544 41
rect 604 37 608 41
rect 1664 37 1668 41
rect 1732 37 1736 41
rect 124 28 128 32
rect 1248 24 1252 28
rect 2788 37 2792 41
rect 2852 37 2856 41
rect 2372 28 2376 32
rect 3444 24 3448 28
rect 3932 240 3936 244
rect 3988 240 3992 244
rect 3932 224 3936 228
rect 17892 232 17896 237
rect 17908 2388 17912 2392
rect 17908 736 17912 740
rect 4080 224 4084 228
rect 3976 149 3980 153
rect 4032 136 4036 140
rect 4032 108 4036 112
rect 3516 24 3520 28
rect 4032 24 4036 28
rect 17908 16 17912 20
rect -12 8 -8 12
rect 28 8 32 12
rect 1152 8 1156 12
rect 1152 -24 1156 -20
rect 2276 8 2280 12
rect 2276 -48 2280 -44
rect 3400 8 3404 12
rect 3400 -72 3404 -68
use 8in-multiplier  8in-multiplier_0
timestamp 1653419601
transform 1 0 15402 0 1 717
box 180 0 2432 280
use 16in-multiplicand  16in-multiplicand_0
timestamp 1653419554
transform 1 0 -181 0 1 2355
box 184 12 4684 292
use 16in-product  16in-product_0
timestamp 1653419529
transform 1 0 2768 0 1 -16
box -2768 16 1712 312
use alu16bit  alu16bit_0
timestamp 1653298574
transform 1 0 4843 0 1 1367
box -8812 -12 8656 224
<< labels >>
rlabel m2contact -102 2520 -98 2524 1 A8
rlabel m2contact -100 2408 -96 2412 1 A0
rlabel m2contact 619 2330 623 2334 1 A1
rlabel m2contact 1211 2344 1215 2348 1 A2
rlabel m2contact 1747 2336 1751 2340 1 A3
rlabel m2contact 2339 2342 2343 2346 1 A4
rlabel m2contact 2875 2339 2879 2343 1 A5
rlabel m2contact 3467 2347 3471 2351 1 A6
rlabel m2contact 4003 2340 4007 2344 1 A7
rlabel m2contact 3956 2700 3960 2704 1 A15
rlabel m2contact 3365 2701 3369 2705 1 A14
rlabel m2contact 2827 2704 2831 2708 1 A13
rlabel m2contact 2239 2700 2243 2704 1 A12
rlabel m2contact 1699 2702 1703 2706 1 A11
rlabel m2contact 1108 2696 1112 2700 1 A10
rlabel m2contact 571 2684 575 2688 1 A9
rlabel m2contact 17278 1036 17282 1040 1 B4
rlabel m2contact 17326 694 17330 698 1 B0
rlabel m2contact 16707 696 16711 700 1 B1
rlabel m2contact 16699 700 16703 704 1 B5
rlabel m2contact 16152 1009 16156 1013 1 B6
rlabel m2contact 16202 695 16206 699 1 B2
rlabel m2contact 15565 757 15569 761 1 B3
rlabel m2contact 15573 870 15577 874 1 B7
rlabel metal1 2312 2667 2316 2671 1 s_0
rlabel metal1 2312 2655 2316 2659 1 reset_0
rlabel metal1 2312 2639 2316 2643 1 phi1_0
rlabel metal1 2312 2619 2316 2623 1 phi2_0
rlabel metal2 4592 2603 4596 2607 1 Vdd
rlabel metal2 4597 2387 4601 2391 1 Gnd
rlabel metal1 17244 993 17248 997 1 s_1
rlabel metal1 17244 985 17248 989 1 reset_1
rlabel metal1 17244 977 17248 981 1 phi1_1
rlabel metal1 17244 969 17248 973 1 phi2_1
rlabel metal1 3912 272 3916 276 1 s_2
rlabel metal1 3912 264 3916 268 1 reset_2
rlabel metal1 3912 256 3916 260 1 phi1_2
rlabel metal1 3912 248 3916 252 1 phi2_2
rlabel metal1 552 186 556 189 1 q15
rlabel metal1 1088 186 1092 189 1 q14
rlabel metal1 1676 186 1680 189 1 q13
rlabel metal1 2212 186 2216 189 1 q12
rlabel metal1 2800 188 2804 191 1 q11
rlabel metal1 3336 188 3340 191 1 q10
rlabel metal1 3924 192 3928 195 1 q9
rlabel metal1 4460 193 4464 196 1 q8
rlabel metal1 4460 55 4464 58 1 q0
rlabel metal1 3924 51 3928 54 1 q1
rlabel metal1 3336 52 3340 55 1 q2
rlabel metal1 2800 61 2804 64 1 q3
rlabel metal1 2212 68 2216 71 1 q4
rlabel metal1 1676 66 1680 69 1 q5
rlabel metal1 1088 61 1092 64 1 q6
rlabel metal1 552 57 556 60 1 q7
<< end >>
