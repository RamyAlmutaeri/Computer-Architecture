magic
tech scmos
timestamp 1652698805
<< polysilicon >>
rect 16 100 18 102
rect 28 100 30 102
rect 16 76 18 96
rect 12 74 18 76
rect 16 12 18 74
rect 28 60 30 96
rect 28 12 30 56
rect 16 6 18 8
rect 28 6 30 8
<< ndiffusion >>
rect 12 8 16 12
rect 18 8 28 12
rect 30 8 32 12
rect 36 8 40 12
<< pdiffusion >>
rect 12 96 16 100
rect 18 96 20 100
rect 24 96 28 100
rect 30 96 36 100
<< metal1 >>
rect 20 100 24 104
rect 8 92 12 96
rect 36 92 40 96
rect 8 88 40 92
rect 36 60 40 88
rect 8 56 28 60
rect 36 56 52 60
rect 64 56 76 60
rect 36 20 40 56
rect 8 16 40 20
rect 8 12 12 16
rect 32 4 36 8
<< metal2 >>
rect 0 104 20 108
rect 24 104 40 108
rect 76 104 84 108
rect 0 0 32 4
rect 36 0 40 4
rect 76 0 84 4
<< ntransistor >>
rect 16 8 18 12
rect 28 8 30 12
<< ptransistor >>
rect 16 96 18 100
rect 28 96 30 100
<< polycontact >>
rect 8 72 12 76
rect 28 56 32 60
<< ndcontact >>
rect 8 8 12 12
rect 32 8 36 12
<< pdcontact >>
rect 8 96 12 100
rect 20 96 24 100
rect 36 96 40 100
<< m2contact >>
rect 20 104 24 108
rect 32 0 36 4
use inverter  inverter_0
timestamp 1652558825
transform 1 0 40 0 1 0
box 0 0 36 108
<< end >>
