magic
tech scmos
timestamp 1653253929
<< polysilicon >>
rect 8 60 10 62
rect 40 60 42 62
rect 8 40 10 56
rect 4 38 10 40
rect 8 12 10 38
rect 40 40 42 56
rect 40 12 42 36
rect 8 6 10 8
rect 40 6 42 8
<< ndiffusion >>
rect 4 8 8 12
rect 10 8 20 12
rect 32 8 40 12
rect 42 8 52 12
<< pdiffusion >>
rect 4 56 8 60
rect 10 56 20 60
rect 32 56 40 60
rect 42 56 52 60
<< metal1 >>
rect 0 60 4 64
rect 28 60 32 64
rect 20 40 24 56
rect 20 36 40 40
rect 20 12 24 36
rect 52 12 56 56
rect 0 4 4 8
rect 28 4 32 8
<< metal2 >>
rect 4 64 28 68
rect 32 64 56 68
rect 4 0 28 4
rect 32 0 56 4
<< ntransistor >>
rect 8 8 10 12
rect 40 8 42 12
<< ptransistor >>
rect 8 56 10 60
rect 40 56 42 60
<< polycontact >>
rect 0 36 4 40
rect 40 36 44 40
<< ndcontact >>
rect 0 8 4 12
rect 20 8 24 12
rect 28 8 32 12
rect 52 8 56 12
<< pdcontact >>
rect 0 56 4 60
rect 20 56 24 60
rect 28 56 32 60
rect 52 56 56 60
<< m2contact >>
rect 0 64 4 68
rect 28 64 32 68
rect 0 0 4 4
rect 28 0 32 4
<< end >>
