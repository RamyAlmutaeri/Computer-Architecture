magic
tech scmos
timestamp 1653295885
<< metal1 >>
rect -384 232 120 236
rect 116 208 120 232
rect -188 200 92 204
rect 140 200 692 204
rect 732 200 908 204
rect 4192 200 4196 204
rect 3996 184 4000 188
rect -3900 100 -3896 104
rect -2816 100 -2812 104
rect -1700 100 -1696 104
rect -616 100 -612 104
rect 484 100 488 104
rect 1568 100 1572 104
rect 2684 100 2688 104
rect 3768 100 3772 104
rect -3376 92 -3372 96
rect -2292 92 -2288 96
rect -1176 92 -1172 96
rect -92 92 -88 96
rect 1008 92 1012 96
rect 2092 92 2096 96
rect 3208 92 3212 96
rect 4292 92 4296 96
rect -3900 76 -3896 80
rect -2816 76 -2812 80
rect -1700 76 -1696 80
rect -616 76 -612 80
rect 484 76 488 80
rect 1568 76 1572 80
rect 2684 76 2688 80
rect 3768 76 3772 80
<< metal2 >>
rect -388 188 -384 232
rect 96 200 136 204
rect 696 200 728 204
rect -92 140 28 144
rect 4288 140 4292 144
rect -92 36 28 40
rect 4288 36 4292 40
<< m2contact >>
rect -388 232 -384 236
rect 92 200 96 204
rect 136 200 140 204
rect 692 200 696 204
rect 728 200 732 204
rect -388 184 -384 188
use nal4bit  nal4bit_0
timestamp 1653255048
transform 1 0 2192 0 1 4
box -2196 0 2104 232
use nal4bit  nal4bit_1
timestamp 1653255048
transform 1 0 -2192 0 1 4
box -2196 0 2104 232
<< end >>
