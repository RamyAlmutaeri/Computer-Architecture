magic
tech scmos
timestamp 1652541516
<< polysilicon >>
rect 16 100 18 102
rect 24 100 26 102
rect 40 100 42 102
rect 48 100 50 102
rect 60 100 62 102
rect 16 60 18 96
rect 24 70 26 96
rect 24 68 34 70
rect 12 58 18 60
rect 16 12 18 58
rect 24 52 26 56
rect 32 51 34 68
rect 40 60 42 96
rect 48 60 50 96
rect 60 84 62 96
rect 32 48 42 51
rect 24 12 26 48
rect 40 44 42 48
rect 40 12 42 40
rect 48 12 50 56
rect 60 28 62 80
rect 60 12 62 24
rect 16 6 18 8
rect 24 6 26 8
rect 40 6 42 8
rect 48 6 50 8
rect 60 6 62 8
<< ndiffusion >>
rect 12 8 16 12
rect 18 8 24 12
rect 26 8 32 12
rect 36 8 40 12
rect 42 8 48 12
rect 50 8 52 12
rect 56 8 60 12
rect 62 8 68 12
<< pdiffusion >>
rect 12 96 16 100
rect 18 96 24 100
rect 26 96 32 100
rect 36 96 40 100
rect 42 96 48 100
rect 50 96 52 100
rect 56 96 60 100
rect 62 96 68 100
<< metal1 >>
rect 8 100 12 104
rect 52 100 56 104
rect 32 84 36 96
rect 32 80 60 84
rect 68 60 72 96
rect 28 56 40 60
rect 52 56 72 60
rect 8 48 24 52
rect 8 40 40 44
rect 32 24 60 28
rect 32 12 36 24
rect 68 12 72 56
rect 8 4 12 8
rect 52 4 56 8
<< metal2 >>
rect 0 104 8 108
rect 12 104 52 108
rect 56 104 80 108
rect 0 0 8 4
rect 12 0 52 4
rect 56 0 80 4
<< ntransistor >>
rect 16 8 18 12
rect 24 8 26 12
rect 40 8 42 12
rect 48 8 50 12
rect 60 8 62 12
<< ptransistor >>
rect 16 96 18 100
rect 24 96 26 100
rect 40 96 42 100
rect 48 96 50 100
rect 60 96 62 100
<< polycontact >>
rect 8 56 12 60
rect 24 56 28 60
rect 24 48 28 52
rect 60 80 64 84
rect 40 56 44 60
rect 48 56 52 60
rect 40 40 44 44
rect 60 24 64 28
<< ndcontact >>
rect 8 8 12 12
rect 32 8 36 12
rect 52 8 56 12
rect 68 8 72 12
<< pdcontact >>
rect 8 96 12 100
rect 32 96 36 100
rect 52 96 56 100
rect 68 96 72 100
<< m2contact >>
rect 8 104 12 108
rect 52 104 56 108
rect 8 0 12 4
rect 52 0 56 4
<< end >>
