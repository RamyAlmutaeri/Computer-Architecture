magic
tech scmos
timestamp 1653419554
<< metal1 >>
rect 760 288 1323 292
rect 1889 288 2452 292
rect 3017 288 3580 292
rect 876 280 1308 284
rect 208 212 224 215
rect 1336 212 1352 215
rect 2464 212 2484 215
rect 3592 212 3612 215
rect 184 16 188 212
rect 744 200 748 212
rect 1280 200 1284 212
rect 1872 200 1876 212
rect 2408 200 2412 212
rect 3000 200 3004 212
rect 3536 200 3540 212
rect 4128 200 4132 212
rect 4664 200 4668 204
rect 264 165 268 169
rect 800 165 804 169
rect 1392 165 1396 169
rect 1928 165 1932 169
rect 2520 165 2524 169
rect 3056 165 3060 169
rect 3648 165 3652 169
rect 4184 165 4188 169
rect 1332 100 1352 103
rect 2460 100 2484 103
rect 3588 100 3604 103
rect 744 88 748 100
rect 1280 88 1284 100
rect 1872 88 1876 100
rect 2408 88 2412 100
rect 3000 88 3004 100
rect 3536 88 3540 100
rect 4128 88 4132 100
rect 264 53 268 57
rect 800 53 804 57
rect 1392 53 1396 57
rect 1928 53 1932 57
rect 2520 53 2524 57
rect 3056 53 3060 57
rect 3648 53 3652 57
rect 4184 53 4188 57
rect 4664 16 4668 92
rect 184 12 4668 16
<< metal2 >>
rect 1312 280 1492 284
rect 2024 280 2620 284
rect 3152 280 3748 284
rect 888 272 1484 276
rect 2016 272 2612 276
rect 3144 272 3740 276
rect 880 264 1472 268
rect 2008 264 2600 268
rect 3136 264 3728 268
rect 1296 248 1348 252
rect 2424 248 2476 252
rect 3552 248 3604 252
rect 188 212 204 215
rect 228 212 264 215
rect 748 212 800 215
rect 1284 212 1332 215
rect 1356 212 1392 215
rect 1876 212 1928 215
rect 2412 212 2460 215
rect 2488 212 2520 215
rect 3004 212 3055 215
rect 3540 212 3588 215
rect 3616 212 3648 215
rect 4132 212 4184 215
rect 1872 211 1932 212
rect 208 99 264 103
rect 748 100 800 103
rect 1284 100 1328 103
rect 1356 100 1392 103
rect 1876 100 1928 103
rect 2412 100 2456 103
rect 2488 100 2520 103
rect 3004 100 3056 103
rect 3540 100 3584 103
rect 3608 100 3648 103
rect 4132 100 4184 103
rect 1296 32 1348 36
rect 2424 32 2476 36
rect 3552 32 3604 36
<< m2contact >>
rect 1308 280 1312 284
rect 2020 280 2024 284
rect 3148 280 3152 284
rect 884 272 888 276
rect 2012 272 2016 276
rect 3140 272 3144 276
rect 876 264 880 268
rect 1472 264 1476 268
rect 2004 264 2008 268
rect 2600 264 2604 268
rect 3132 264 3136 268
rect 3728 264 3732 268
rect 184 212 188 216
rect 204 212 208 216
rect 224 212 228 216
rect 264 212 268 216
rect 744 212 748 216
rect 800 212 804 216
rect 1280 212 1284 216
rect 1332 212 1336 216
rect 1352 212 1356 216
rect 1392 212 1396 216
rect 1872 212 1876 216
rect 1928 212 1932 216
rect 2408 212 2412 216
rect 2460 212 2464 216
rect 2484 212 2488 216
rect 2520 212 2524 216
rect 3000 212 3004 216
rect 3055 212 3059 216
rect 3536 212 3540 216
rect 3588 212 3592 216
rect 3612 212 3616 216
rect 3648 212 3652 216
rect 4128 212 4132 216
rect 4184 212 4188 216
rect 264 99 268 103
rect 744 100 748 104
rect 800 100 804 104
rect 1280 100 1284 104
rect 1328 100 1332 104
rect 1352 100 1356 104
rect 1392 100 1396 104
rect 1872 100 1876 104
rect 1928 100 1932 104
rect 2408 100 2412 104
rect 2456 100 2460 104
rect 2484 100 2488 104
rect 2520 100 2524 104
rect 3000 100 3004 104
rect 3056 100 3060 104
rect 3536 100 3540 104
rect 3584 100 3588 104
rect 3604 100 3608 104
rect 3648 100 3652 104
rect 4128 100 4132 104
rect 4184 100 4188 104
use 4in-multiplicand  4in-multiplicand_0
timestamp 1653191793
transform 1 0 900 0 1 144
box -708 -120 400 148
use 4in-multiplicand  4in-multiplicand_1
timestamp 1653191793
transform 1 0 2028 0 1 144
box -708 -120 400 148
use 4in-multiplicand  4in-multiplicand_2
timestamp 1653191793
transform 1 0 3156 0 1 144
box -708 -120 400 148
use 4in-multiplicand  4in-multiplicand_3
timestamp 1653191793
transform 1 0 4284 0 1 144
box -708 -120 400 148
<< end >>
