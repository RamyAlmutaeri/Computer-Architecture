magic
tech scmos
timestamp 1652779389
<< polysilicon >>
rect 16 92 19 94
rect 16 12 19 88
rect 16 5 19 8
<< ndiffusion >>
rect 8 8 16 12
rect 19 8 36 12
rect 40 8 52 12
<< pdiffusion >>
rect 8 88 16 92
rect 19 88 36 92
rect 40 88 52 92
<< metal1 >>
rect 4 92 8 96
rect 36 12 40 88
rect 4 4 8 8
<< metal2 >>
rect 0 96 4 100
rect 8 96 56 100
rect 0 0 4 4
rect 8 0 56 4
<< ntransistor >>
rect 16 8 19 12
<< ptransistor >>
rect 16 88 19 92
<< ndcontact >>
rect 4 8 8 12
rect 36 8 40 12
<< pdcontact >>
rect 4 88 8 92
rect 36 88 40 92
<< m2contact >>
rect 4 96 8 100
rect 4 0 8 4
<< end >>
