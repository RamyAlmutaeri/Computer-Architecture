magic
tech scmos
timestamp 1653250592
<< metal1 >>
rect -4 200 124 204
rect -196 196 -20 200
rect -4 192 0 200
rect 140 196 696 200
rect 744 196 916 200
rect 2000 196 2004 200
rect -276 188 -216 192
rect -180 188 0 192
rect -276 184 -272 188
rect -392 180 -272 184
rect 1804 180 1808 184
rect -1708 96 -1704 100
rect -624 96 -620 100
rect 492 96 496 100
rect 1576 96 1580 100
rect -1184 88 -1180 92
rect -100 88 -96 92
rect 1016 88 1020 92
rect 2100 88 2104 92
rect -1708 72 -1704 76
rect -624 72 -620 76
rect 492 72 496 76
rect 1576 72 1580 76
<< metal2 >>
rect -16 196 136 200
rect 700 196 740 200
rect -212 188 -184 192
rect -100 136 36 140
rect 2096 136 2100 140
rect -100 32 36 36
rect 2096 32 2100 36
<< m2contact >>
rect -20 196 -16 200
rect 136 196 140 200
rect 696 196 700 200
rect 740 196 744 200
rect -216 188 -212 192
rect -184 188 -180 192
use nalu2bit  nalu2bit_0
timestamp 1653247424
transform 1 0 1088 0 1 0
box -1084 0 1016 232
use nalu2bit  nalu2bit_1
timestamp 1653247424
transform 1 0 -1112 0 1 0
box -1084 0 1016 232
<< labels >>
rlabel metal1 2000 196 2004 200 1 E
rlabel metal1 1804 180 1808 184 1 Cin
rlabel metal1 1576 96 1580 100 1 A0
rlabel metal1 1016 88 1020 92 1 D1
rlabel metal1 -100 88 -96 92 1 D2
rlabel metal1 -1184 88 -1180 92 1 D3
rlabel metal1 492 96 496 100 1 A1
rlabel metal1 492 72 496 76 1 B1
rlabel metal1 -624 96 -620 100 1 A2
rlabel metal1 -624 72 -620 76 1 B2
rlabel metal1 -1708 96 -1704 100 1 A3
rlabel metal1 -1708 72 -1704 76 1 B3
rlabel metal2 2096 136 2100 140 1 Vdd
rlabel metal2 2096 32 2100 36 1 Gnd
rlabel metal1 1576 72 1580 76 1 B0
rlabel metal1 2100 88 2104 92 7 D0
<< end >>
