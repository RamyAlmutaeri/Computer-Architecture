magic
tech scmos
timestamp 1653419779
<< metal1 >>
rect -528 162 -524 516
rect -516 98 -512 528
rect -504 154 -500 540
rect -504 4 -500 150
rect -492 106 -488 552
rect -492 -48 -488 102
rect -480 146 -476 564
rect -480 -4 -476 142
rect -480 -151 -476 -8
rect -468 114 -464 576
rect -468 -32 -464 110
rect -468 -175 -464 -36
rect -456 138 -452 588
rect -456 -24 -452 134
rect -456 -167 -452 -28
rect -444 122 -440 600
rect -107 499 -101 501
rect -107 495 -106 499
rect -102 495 -101 499
rect 488 499 492 508
rect -204 381 -199 432
rect -118 395 -112 397
rect -118 391 -117 395
rect -113 391 -112 395
rect -118 280 -112 391
rect -118 276 -117 280
rect -113 276 -112 280
rect -308 158 -303 162
rect -118 161 -112 276
rect -444 -40 -440 118
rect -118 157 -117 161
rect -113 157 -112 161
rect -118 64 -112 157
rect -118 60 -117 64
rect -113 60 -112 64
rect -118 42 -112 60
rect -118 38 -117 42
rect -113 38 -112 42
rect -302 0 -296 4
rect -300 -8 -297 -4
rect -143 -12 -125 -8
rect -300 -28 -297 -24
rect -300 -36 -298 -32
rect -300 -44 -297 -40
rect -444 -127 -440 -44
rect -300 -52 -297 -48
rect -118 -85 -112 38
rect -118 -89 -117 -85
rect -113 -89 -112 -85
rect -444 -224 -440 -131
rect -118 -135 -112 -89
rect -107 384 -101 495
rect 614 491 618 508
rect 753 499 757 516
rect 76 483 84 484
rect 76 479 78 483
rect 83 479 84 483
rect -107 380 -106 384
rect -102 380 -101 384
rect -107 265 -101 380
rect -107 261 -106 265
rect -102 261 -101 265
rect -107 182 -101 261
rect -107 178 -106 182
rect -102 178 -101 182
rect -107 146 -101 178
rect -107 142 -106 146
rect -102 142 -101 146
rect -107 32 -101 142
rect -107 28 -106 32
rect -102 28 -101 32
rect -107 5 -101 28
rect -107 1 -106 5
rect -102 1 -101 5
rect -107 -95 -101 1
rect -52 130 -48 455
rect 65 447 71 448
rect 65 443 66 447
rect 70 443 71 447
rect 65 437 71 443
rect 65 432 66 437
rect 70 432 71 437
rect 49 427 55 429
rect 49 423 50 427
rect 54 423 55 427
rect -52 -59 -48 126
rect -40 -67 -36 340
rect 49 312 55 423
rect 49 308 50 312
rect 54 308 55 312
rect 49 256 55 308
rect 49 252 50 256
rect 54 252 55 256
rect -107 -99 -106 -95
rect -102 -99 -101 -95
rect -107 -100 -101 -99
rect -30 -75 -26 221
rect 49 193 55 252
rect 49 189 50 193
rect 54 189 55 193
rect -30 -119 -26 -79
rect -17 -51 -13 102
rect 49 74 55 189
rect 65 328 71 432
rect 65 324 66 328
rect 70 324 71 328
rect 65 209 71 324
rect 65 205 66 209
rect 70 205 71 209
rect 65 93 71 205
rect 76 368 84 479
rect 76 364 78 368
rect 83 364 84 368
rect 76 249 84 364
rect 76 245 78 249
rect 83 245 84 249
rect 76 131 84 245
rect 76 126 78 131
rect 82 126 84 131
rect 76 125 84 126
rect 510 480 515 487
rect 510 476 532 480
rect 510 459 515 476
rect 615 455 626 459
rect 510 360 515 455
rect 764 443 768 528
rect 622 417 626 429
rect 523 395 527 404
rect 612 387 616 391
rect 600 369 605 379
rect 510 351 515 356
rect 510 347 529 351
rect 510 243 515 347
rect 616 346 620 356
rect 616 342 629 346
rect 625 336 629 342
rect 776 336 780 540
rect 788 321 792 552
rect 600 265 605 275
rect 510 234 515 239
rect 510 230 523 234
rect 510 126 515 230
rect 608 228 612 239
rect 608 224 621 228
rect 617 219 621 224
rect 800 218 804 564
rect 812 203 816 576
rect 510 116 515 122
rect 510 112 526 116
rect 608 112 612 122
rect 608 108 620 112
rect 616 101 620 108
rect 824 100 828 588
rect 65 89 66 93
rect 70 89 71 93
rect 65 88 71 89
rect 836 88 840 600
rect 49 70 50 74
rect 54 70 55 74
rect 49 68 55 70
rect 616 65 620 74
rect -17 -54 98 -51
rect -17 -55 78 -54
rect 87 -55 98 -54
rect -118 -139 -117 -135
rect -113 -139 -112 -135
rect -118 -199 -112 -139
rect -17 -224 -13 -55
rect 6 -63 7 -59
rect 11 -63 94 -59
rect 205 -64 213 -59
rect -4 -71 94 -67
<< metal2 >>
rect -440 600 836 604
rect -452 588 824 592
rect -464 576 812 580
rect -476 564 800 568
rect -488 552 788 556
rect -500 540 776 544
rect -512 528 764 532
rect -524 516 753 520
rect 492 508 526 512
rect 603 508 614 512
rect -102 495 85 499
rect 591 495 753 499
rect 83 479 100 483
rect -48 455 104 459
rect 515 455 611 459
rect 491 447 531 451
rect 70 443 100 447
rect 100 439 101 443
rect 691 439 764 443
rect -199 432 66 437
rect 54 423 101 427
rect 436 413 622 417
rect -113 391 88 395
rect 491 391 523 395
rect 527 391 612 395
rect -102 380 84 384
rect 488 379 521 383
rect 83 364 100 368
rect 605 365 633 369
rect 515 356 616 360
rect -36 340 103 344
rect 487 332 529 336
rect 599 332 776 336
rect 70 324 100 328
rect 695 317 788 321
rect 54 308 100 312
rect 625 302 629 305
rect 488 298 629 302
rect -113 276 85 280
rect 488 275 521 279
rect -102 261 84 265
rect 487 261 513 265
rect -212 252 50 256
rect 591 251 596 266
rect 605 261 633 265
rect 83 245 99 249
rect 591 247 609 251
rect 515 239 608 243
rect -26 221 104 225
rect 491 213 519 217
rect 588 214 800 218
rect 70 205 100 209
rect 684 199 812 203
rect 54 189 100 193
rect 500 187 616 191
rect 500 184 505 187
rect -132 178 -106 182
rect 490 180 505 184
rect -524 158 -312 162
rect -113 157 83 161
rect 489 157 515 161
rect 586 158 612 162
rect -500 150 -304 154
rect -476 142 -304 146
rect -102 142 84 146
rect 490 142 521 146
rect -452 134 -304 138
rect 598 135 602 147
rect 607 143 612 158
rect 598 131 614 135
rect -144 126 -52 130
rect 82 126 99 130
rect 515 122 608 126
rect -440 118 -302 122
rect -464 110 -303 114
rect -488 102 -303 106
rect -13 102 104 106
rect -512 94 -304 98
rect 489 94 526 98
rect 595 96 824 100
rect 70 89 101 92
rect 685 83 836 87
rect 54 70 99 74
rect -132 60 -117 64
rect 491 61 616 64
rect -113 38 82 42
rect 489 38 523 42
rect 600 32 604 44
rect -135 28 -106 32
rect 600 28 614 32
rect -500 0 -306 4
rect -102 1 98 5
rect -476 -8 -304 -4
rect -121 -12 -44 -8
rect 94 -15 98 1
rect -452 -28 -304 -24
rect -464 -36 -304 -32
rect -440 -44 -304 -40
rect -488 -52 -304 -48
rect -48 -63 7 -59
rect -36 -71 -8 -67
rect -26 -79 91 -75
rect -134 -89 -117 -85
rect -216 -99 -106 -95
rect -258 -124 -30 -119
rect -440 -131 -294 -127
rect 94 -135 98 -115
rect -113 -139 98 -135
rect -476 -155 -294 -151
rect -452 -171 -294 -167
rect -464 -179 -290 -175
rect -217 -203 -118 -199
rect -440 -228 -17 -224
<< m2contact >>
rect -444 600 -440 604
rect -456 588 -452 592
rect -468 576 -464 580
rect -480 564 -476 568
rect -492 552 -488 556
rect -504 540 -500 544
rect -516 528 -512 532
rect -528 516 -524 520
rect -528 158 -524 162
rect -516 94 -512 98
rect -504 150 -500 154
rect -504 0 -500 4
rect -492 102 -488 106
rect -492 -52 -488 -48
rect -480 142 -476 146
rect -480 -8 -476 -4
rect -480 -155 -476 -151
rect -468 110 -464 114
rect -468 -36 -464 -32
rect -456 134 -452 138
rect -456 -28 -452 -24
rect -456 -171 -452 -167
rect 836 600 840 604
rect 824 588 828 592
rect 812 576 816 580
rect 800 564 804 568
rect 788 552 792 556
rect 776 540 780 544
rect 764 528 768 532
rect 753 516 757 520
rect 488 508 492 512
rect -106 495 -102 499
rect 614 508 618 512
rect 488 495 492 499
rect 587 495 591 499
rect -204 432 -199 437
rect -117 391 -113 395
rect -117 276 -113 280
rect -312 158 -308 162
rect -444 118 -440 122
rect -117 157 -113 161
rect -117 60 -113 64
rect -117 38 -113 42
rect -306 0 -302 4
rect -304 -8 -300 -4
rect -125 -12 -121 -8
rect -304 -28 -300 -24
rect -304 -36 -300 -32
rect -444 -44 -440 -40
rect -304 -44 -300 -40
rect -304 -52 -300 -48
rect -117 -89 -113 -85
rect -444 -131 -440 -127
rect -294 -131 -290 -127
rect -468 -179 -464 -175
rect 753 495 757 499
rect 614 487 618 491
rect 78 479 83 483
rect -106 380 -102 384
rect -106 261 -102 265
rect -106 178 -102 182
rect -106 142 -102 146
rect -106 28 -102 32
rect -106 1 -102 5
rect -52 455 -48 459
rect 66 443 70 447
rect 66 432 70 437
rect 50 423 54 427
rect -52 126 -48 130
rect -40 340 -36 344
rect -44 -12 -40 -8
rect -52 -63 -48 -59
rect 50 308 54 312
rect 50 252 54 256
rect -40 -71 -36 -67
rect -30 221 -26 225
rect -106 -99 -102 -95
rect 50 189 54 193
rect -30 -79 -26 -75
rect -30 -124 -26 -119
rect -17 102 -13 106
rect 66 324 70 328
rect 66 205 70 209
rect 78 364 83 368
rect 78 245 83 249
rect 78 126 82 131
rect 510 455 515 459
rect 611 455 615 459
rect 531 447 535 451
rect 687 439 691 443
rect 764 439 768 443
rect 622 413 626 417
rect 523 404 527 408
rect 523 391 527 395
rect 612 391 616 395
rect 612 383 616 387
rect 600 379 605 383
rect 600 365 605 369
rect 510 356 515 360
rect 616 356 620 360
rect 529 332 533 336
rect 594 331 599 336
rect 776 332 780 336
rect 690 317 695 321
rect 788 317 792 321
rect 625 305 629 309
rect 600 275 605 279
rect 600 261 605 265
rect 510 239 515 243
rect 608 239 612 243
rect 519 213 523 217
rect 584 214 588 218
rect 800 214 804 218
rect 680 199 684 203
rect 812 199 816 203
rect 616 187 621 191
rect 510 122 515 126
rect 608 122 612 126
rect 526 94 530 98
rect 590 96 595 100
rect 824 96 828 100
rect 66 89 70 93
rect 680 83 685 87
rect 836 83 840 88
rect 50 70 54 74
rect 616 61 620 65
rect -117 -139 -113 -135
rect -294 -155 -290 -151
rect -294 -171 -290 -167
rect -118 -203 -112 -199
rect -444 -228 -440 -224
rect 7 -63 11 -59
rect -8 -71 -4 -67
rect 91 -79 95 -75
rect -17 -228 -13 -224
use 2inAND  2inAND_0
timestamp 1653329418
transform 1 0 523 0 1 404
box 0 0 84 108
use 2inAND  2inAND_1
timestamp 1653329418
transform 1 0 614 0 1 383
box 0 0 84 108
use 2inAND  2inAND_2
timestamp 1653329418
transform 1 0 521 0 1 275
box 0 0 84 108
use 2inAND  2inAND_3
timestamp 1653329418
transform 1 0 617 0 1 261
box 0 0 84 108
use 2inAND  2inAND_4
timestamp 1653329418
transform 1 0 511 0 1 158
box 0 0 84 108
use 2inAND  2inAND_5
timestamp 1653329418
transform 1 0 609 0 1 143
box 0 0 84 108
use 2inAND  2inAND_6
timestamp 1653329418
transform 1 0 518 0 1 40
box 0 0 84 108
use 2inAND  2inAND_7
timestamp 1653329418
transform 1 0 608 0 1 27
box 0 0 84 108
use 4inAND  4inAND_1
timestamp 1653262109
transform 1 0 94 0 1 -119
box 0 0 112 108
use dflipflopER  dflipflopER_0
timestamp 1653329719
transform 1 0 -74 0 1 38
box 156 0 565 108
use dflipflopER  dflipflopER_1
timestamp 1653329719
transform 1 0 -73 0 1 157
box 156 0 565 108
use dflipflopER  dflipflopER_2
timestamp 1653329719
transform 1 0 -73 0 1 276
box 156 0 565 108
use dflipflopER  dflipflopER_3
timestamp 1653329719
transform 1 0 -72 0 1 391
box 156 0 565 108
use nxta  nxta_0
timestamp 1653244860
transform 1 0 -290 0 1 60
box -15 0 158 122
use nxtb  nxtb_0
timestamp 1653204617
transform 1 0 -290 0 1 -80
box -16 -9 156 112
use xnor  xnor_0
timestamp 1652719145
transform 1 0 -282 0 1 -195
box -16 -8 68 100
<< labels >>
rlabel metal1 88 -53 88 -53 1 nxtd
rlabel metal1 208 -62 208 -62 1 nextEn
rlabel metal1 90 -61 90 -61 1 nxta
rlabel metal1 90 -69 90 -69 1 nxtb
rlabel m2contact 92 -77 92 -77 1 nxtc
rlabel metal1 -202 383 -202 383 1 phi1
rlabel metal2 -209 254 -209 254 1 phi2
rlabel metal1 512 485 512 485 1 En
rlabel m2contact -114 -201 -114 -201 1 gnd
rlabel metal1 -104 -92 -104 -92 1 vdd
rlabel metal1 80 133 80 133 1 reset
<< end >>
