magic
tech scmos
timestamp 1652558825
<< polysilicon >>
rect 16 100 18 102
rect 16 60 18 96
rect 12 58 18 60
rect 16 12 18 58
rect 16 6 18 8
<< ndiffusion >>
rect 12 8 16 12
rect 18 8 24 12
<< pdiffusion >>
rect 12 96 16 100
rect 18 96 24 100
<< metal1 >>
rect 8 100 12 104
rect 24 12 28 96
rect 8 4 12 8
<< metal2 >>
rect 0 104 8 108
rect 12 104 36 108
rect 0 0 8 4
rect 12 0 36 4
<< ntransistor >>
rect 16 8 18 12
<< ptransistor >>
rect 16 96 18 100
<< polycontact >>
rect 8 56 12 60
<< ndcontact >>
rect 8 8 12 12
rect 24 8 28 12
<< pdcontact >>
rect 8 96 12 100
rect 24 96 28 100
<< m2contact >>
rect 8 104 12 108
rect 8 0 12 4
<< end >>
