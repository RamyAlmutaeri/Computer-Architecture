magic
tech scmos
timestamp 1653418476
<< polysilicon >>
rect 16 100 19 102
rect 16 12 19 96
rect 16 5 19 8
<< ndiffusion >>
rect 8 8 16 12
rect 19 8 36 12
rect 40 8 52 12
<< pdiffusion >>
rect 8 96 16 100
rect 19 96 36 100
rect 40 96 52 100
<< metal1 >>
rect 4 100 8 104
rect 36 12 40 96
rect 4 4 8 8
<< metal2 >>
rect 0 104 4 108
rect 8 104 56 108
rect 0 0 4 4
rect 8 0 56 4
<< ntransistor >>
rect 16 8 19 12
<< ptransistor >>
rect 16 96 19 100
<< ndcontact >>
rect 4 8 8 12
rect 36 8 40 12
<< pdcontact >>
rect 4 96 8 100
rect 36 96 40 100
<< m2contact >>
rect 4 104 8 108
rect 4 0 8 4
<< end >>
