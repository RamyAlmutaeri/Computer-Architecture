magic
tech scmos
timestamp 1653422444
<< polysilicon >>
rect 7 114 9 116
rect 35 114 37 116
rect 51 114 53 116
rect 67 114 69 116
rect 82 114 84 116
rect 99 114 101 116
rect 115 114 117 116
rect 139 114 141 116
rect 7 100 9 110
rect -10 98 9 100
rect 7 12 9 98
rect 35 94 37 110
rect 35 12 37 90
rect 51 86 53 110
rect 51 12 53 82
rect 67 78 69 110
rect 67 12 69 74
rect 82 62 84 110
rect 82 12 84 58
rect 99 54 101 110
rect 99 12 101 50
rect 115 46 117 110
rect 115 12 117 42
rect 139 38 141 110
rect 139 12 141 34
rect 7 6 9 8
rect 35 6 37 8
rect 51 6 53 8
rect 67 6 69 8
rect 82 6 84 8
rect 99 6 101 8
rect 115 6 117 8
rect 139 6 141 8
<< ndiffusion >>
rect -11 8 -1 12
rect 3 8 7 12
rect 9 8 12 12
rect 16 8 18 12
rect 26 8 28 12
rect 32 8 35 12
rect 37 8 42 12
rect 46 8 51 12
rect 53 8 58 12
rect 62 8 67 12
rect 69 8 74 12
rect 78 8 82 12
rect 84 8 99 12
rect 101 8 115 12
rect 117 8 120 12
rect 124 8 126 12
rect 131 8 133 12
rect 137 8 139 12
rect 141 8 146 12
rect 150 8 154 12
<< pdiffusion >>
rect -11 110 -1 114
rect 3 110 7 114
rect 9 110 35 114
rect 37 110 51 114
rect 53 110 67 114
rect 69 110 74 114
rect 78 110 82 114
rect 84 110 90 114
rect 94 110 99 114
rect 101 110 106 114
rect 110 110 115 114
rect 117 110 122 114
rect 126 110 139 114
rect 141 110 146 114
rect 150 110 154 114
<< metal1 >>
rect 74 114 78 118
rect 106 114 110 118
rect -1 70 3 110
rect 90 106 94 110
rect 122 106 126 110
rect 32 90 34 94
rect 48 82 50 86
rect 64 74 66 78
rect -1 12 3 66
rect 146 70 150 110
rect 76 58 80 62
rect 92 50 97 54
rect 108 42 113 46
rect 132 34 137 38
rect 12 12 16 16
rect 28 12 32 24
rect 58 12 62 24
rect 120 12 124 16
rect 133 12 137 24
rect 146 12 150 66
rect 42 4 46 8
rect 74 4 78 8
<< metal2 >>
rect -15 118 74 122
rect 78 118 106 122
rect 110 118 158 122
rect 94 102 122 106
rect -14 90 28 94
rect -14 82 44 86
rect -14 74 60 78
rect -4 66 -1 70
rect 3 66 146 70
rect 150 66 154 70
rect -14 58 72 62
rect -14 50 88 54
rect -14 42 104 46
rect -14 34 128 38
rect 32 24 58 28
rect 62 24 133 28
rect 16 16 120 20
rect -15 0 42 4
rect 46 0 74 4
rect 78 0 158 4
<< ntransistor >>
rect 7 8 9 12
rect 35 8 37 12
rect 51 8 53 12
rect 67 8 69 12
rect 82 8 84 12
rect 99 8 101 12
rect 115 8 117 12
rect 139 8 141 12
<< ptransistor >>
rect 7 110 9 114
rect 35 110 37 114
rect 51 110 53 114
rect 67 110 69 114
rect 82 110 84 114
rect 99 110 101 114
rect 115 110 117 114
rect 139 110 141 114
<< polycontact >>
rect -14 98 -10 102
rect 34 90 38 94
rect 50 82 54 86
rect 66 74 70 78
rect 80 58 84 62
rect 97 50 101 54
rect 113 42 117 46
rect 137 34 141 38
<< ndcontact >>
rect -1 8 3 12
rect 12 8 16 12
rect 28 8 32 12
rect 42 8 46 12
rect 58 8 62 12
rect 74 8 78 12
rect 120 8 124 12
rect 133 8 137 12
rect 146 8 150 12
<< pdcontact >>
rect -1 110 3 114
rect 74 110 78 114
rect 90 110 94 114
rect 106 110 110 114
rect 122 110 126 114
rect 146 110 150 114
<< m2contact >>
rect 74 118 78 122
rect 106 118 110 122
rect 90 102 94 106
rect 122 102 126 106
rect 28 90 32 94
rect 44 82 48 86
rect 60 74 64 78
rect -1 66 3 70
rect 146 66 150 70
rect 72 58 76 62
rect 88 50 92 54
rect 104 42 108 46
rect 128 34 132 38
rect 28 24 32 28
rect 12 16 16 20
rect 58 24 62 28
rect 133 24 137 28
rect 120 16 124 20
rect 42 0 46 4
rect 74 0 78 4
<< end >>
