magic
tech scmos
timestamp 1653422461
<< polysilicon >>
rect 12 104 14 106
rect 40 104 42 106
rect 56 104 58 106
rect 86 104 88 106
rect 102 104 104 106
rect 134 104 136 106
rect 12 83 14 100
rect -3 80 14 83
rect 12 3 14 80
rect 40 76 42 100
rect 40 3 42 72
rect 56 56 58 100
rect 56 3 58 52
rect 86 48 88 100
rect 86 3 88 44
rect 102 40 104 100
rect 102 3 104 36
rect 134 32 136 100
rect 134 3 136 28
rect 12 -3 14 -1
rect 40 -3 42 -1
rect 56 -3 58 -1
rect 86 -3 88 -1
rect 102 -3 104 -1
rect 134 -3 136 -1
<< ndiffusion >>
rect -8 -1 3 3
rect 7 -1 12 3
rect 14 -1 19 3
rect 23 -1 26 3
rect 31 -1 34 3
rect 38 -1 40 3
rect 42 -1 48 3
rect 52 -1 56 3
rect 58 -1 60 3
rect 64 -1 68 3
rect 74 -1 80 3
rect 84 -1 86 3
rect 88 -1 102 3
rect 104 -1 108 3
rect 112 -1 117 3
rect 121 -1 124 3
rect 128 -1 134 3
rect 136 -1 145 3
rect 149 -1 152 3
<< pdiffusion >>
rect -8 100 6 104
rect 10 100 12 104
rect 14 100 40 104
rect 42 100 56 104
rect 58 100 60 104
rect 64 100 68 104
rect 76 100 80 104
rect 84 100 86 104
rect 88 100 92 104
rect 96 100 102 104
rect 104 100 108 104
rect 112 100 134 104
rect 136 100 147 104
rect 151 100 152 104
<< metal1 >>
rect 60 104 64 108
rect 92 104 96 108
rect -7 72 -4 76
rect 6 64 10 100
rect 80 96 84 100
rect 108 96 112 100
rect 36 72 39 76
rect 147 64 151 100
rect -8 52 -4 56
rect -8 44 -4 48
rect -8 36 -4 40
rect -8 28 -4 32
rect 3 3 7 60
rect 52 52 54 56
rect 80 44 84 48
rect 96 36 100 40
rect 128 28 132 32
rect 19 3 23 7
rect 34 3 38 15
rect 60 3 64 15
rect 80 3 84 7
rect 124 3 128 15
rect 145 3 149 60
rect 48 -5 52 -1
rect 108 -5 112 -1
<< metal2 >>
rect -16 108 60 112
rect 64 108 92 112
rect 96 108 156 112
rect 84 92 108 96
rect 0 72 32 76
rect 2 60 3 64
rect 10 60 145 64
rect 0 52 48 56
rect 0 44 76 48
rect 0 36 92 40
rect 0 28 124 32
rect 38 15 60 19
rect 64 15 124 19
rect 23 7 80 11
rect -16 -9 48 -5
rect 52 -9 108 -5
rect 112 -9 156 -5
<< ntransistor >>
rect 12 -1 14 3
rect 40 -1 42 3
rect 56 -1 58 3
rect 86 -1 88 3
rect 102 -1 104 3
rect 134 -1 136 3
<< ptransistor >>
rect 12 100 14 104
rect 40 100 42 104
rect 56 100 58 104
rect 86 100 88 104
rect 102 100 104 104
rect 134 100 136 104
<< polycontact >>
rect -7 80 -3 84
rect 39 72 43 76
rect 54 52 58 56
rect 84 44 88 48
rect 100 36 104 40
rect 132 28 136 32
<< ndcontact >>
rect 3 -1 7 3
rect 19 -1 23 3
rect 34 -1 38 3
rect 48 -1 52 3
rect 60 -1 64 3
rect 80 -1 84 3
rect 108 -1 112 3
rect 124 -1 128 3
rect 145 -1 149 3
<< pdcontact >>
rect 6 100 10 104
rect 60 100 64 104
rect 80 100 84 104
rect 92 100 96 104
rect 108 100 112 104
rect 147 100 151 104
<< m2contact >>
rect 60 108 64 112
rect 92 108 96 112
rect -4 72 0 76
rect 80 92 84 96
rect 108 92 112 96
rect 32 72 36 76
rect 3 60 10 64
rect 145 60 151 64
rect -4 52 0 56
rect -4 44 0 48
rect -4 36 0 40
rect -4 28 0 32
rect 48 52 52 56
rect 76 44 80 48
rect 92 36 96 40
rect 124 28 128 32
rect 34 15 38 19
rect 19 7 23 11
rect 60 15 64 19
rect 124 15 128 19
rect 80 7 84 11
rect 48 -9 52 -5
rect 108 -9 112 -5
<< end >>
