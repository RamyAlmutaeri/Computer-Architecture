magic
tech scmos
timestamp 1653423552
<< metal1 >>
rect 311 902 319 904
rect 311 898 314 902
rect 318 898 319 902
rect 311 666 319 898
rect 311 662 313 666
rect 317 662 319 666
rect 311 660 319 662
rect 332 889 340 891
rect 332 885 336 889
rect 332 484 340 885
rect 410 874 416 876
rect 410 870 411 874
rect 415 870 416 874
rect 410 623 416 870
rect 421 858 427 860
rect 421 854 422 858
rect 421 723 427 854
rect 604 842 612 844
rect 604 838 606 842
rect 610 838 612 842
rect 604 706 612 838
rect 1038 708 1043 908
rect 1808 652 1812 898
rect 332 480 333 484
rect 338 480 340 484
rect 332 478 340 480
rect 1820 485 1824 885
rect 1928 874 1932 876
rect 1920 728 1924 854
rect 1928 624 1932 870
rect 2090 712 2094 838
rect 2522 705 2526 716
rect 1038 251 1044 341
rect 736 247 1044 251
rect 2504 340 2527 344
rect 736 197 740 247
rect 877 220 880 247
rect 859 217 880 220
rect 888 202 899 206
rect 736 193 760 197
rect 888 192 892 202
rect 832 184 843 188
rect 964 181 968 190
rect 609 176 612 180
rect 827 177 856 181
rect 2092 178 2096 181
rect 609 167 612 171
rect 739 165 763 169
rect 609 155 612 157
rect 1392 -16 1396 176
rect 2102 174 2103 177
rect 2093 168 2097 171
rect 2224 165 2228 170
rect 2092 156 2096 159
rect 2504 -16 2508 340
<< metal2 >>
rect 319 902 1764 904
rect 318 898 1808 902
rect 319 896 1764 898
rect 340 885 1820 889
rect 415 870 1928 874
rect 427 859 1916 860
rect 422 858 1916 859
rect 427 854 1920 858
rect 1924 854 1925 858
rect 422 852 1916 854
rect 610 838 2090 842
rect 311 662 313 664
rect 317 662 325 664
rect 311 660 325 662
rect 710 225 751 229
rect 832 225 836 236
rect 868 234 892 238
rect 710 213 714 225
rect 863 188 888 192
rect 860 176 899 181
rect 968 176 1392 181
rect 602 147 605 149
rect 2093 148 2097 151
rect 751 113 755 125
rect 832 121 836 132
rect 868 130 891 134
rect 713 109 755 113
rect 1396 -20 2504 -16
<< m2contact >>
rect 314 898 318 902
rect 313 662 317 666
rect 336 885 340 889
rect 411 870 415 874
rect 422 854 427 858
rect 606 838 610 842
rect 1808 898 1812 902
rect 1820 885 1824 889
rect 333 480 338 484
rect 1928 870 1932 874
rect 1920 854 1924 858
rect 1920 724 1924 728
rect 2090 838 2094 842
rect 1928 620 1932 624
rect 1820 479 1824 485
rect 859 188 863 192
rect 888 188 892 192
rect 856 176 860 181
rect 899 176 903 181
rect 964 176 968 181
rect 1392 176 1396 181
rect 1392 -20 1396 -16
rect 2504 -20 2508 -16
use 2inAND  2inAND_0
timestamp 1653422366
transform 1 0 751 0 1 121
box 0 0 84 108
use 2inAND  2inAND_1
timestamp 1653422366
transform 1 0 891 0 1 130
box 0 0 84 108
use dnctr16  dnctr16_0
timestamp 1653419779
transform 1 0 528 0 1 228
box -528 -228 840 604
use dnctr16  dnctr16_1
timestamp 1653419779
transform 1 0 2012 0 1 229
box -528 -228 840 604
use inverter  inverter_0
timestamp 1652558825
transform 1 0 835 0 1 128
box 0 0 36 108
<< labels >>
rlabel metal1 2226 168 2226 168 1 dncounting
rlabel m2contact 858 179 858 179 1 nxtEn
rlabel metal1 834 186 834 186 1 ctrholder
rlabel metal1 336 888 336 888 5 phi2
rlabel metal1 315 894 315 894 5 phi1
rlabel m2contact 413 871 413 871 5 gnd
rlabel m2contact 424 856 424 856 1 vdd
rlabel metal1 608 835 608 835 5 reset
rlabel metal1 2092 156 2096 159 1 d6
rlabel metal2 2093 148 2097 151 1 d5
rlabel metal1 2092 178 2096 181 1 d4
rlabel metal1 609 169 612 171 1 d3
rlabel metal1 609 155 612 157 1 d2
rlabel metal1 609 178 612 180 1 d0
rlabel metal2 602 147 605 149 1 d1
rlabel metal1 2093 168 2097 171 1 d7
<< end >>
